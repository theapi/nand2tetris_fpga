
/**
 * Just a dummy module.
 */
module boolean_arithmatic(out, in);

output out;
input in;

assign out = in;

endmodule
